/*
 * Copyright (c) 2021 Robert Drehmel
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
interface mmr_readwrite_interface#(
	parameter int NREGS
);

localparam int INDEX_WIDTH = $clog2(NREGS);

logic store;
logic [INDEX_WIDTH-1:0] store_idx;
logic [31:0] store_data;
logic [31:0] data [NREGS];

modport master(
	output store,
	output store_idx,
	output store_data,
	input data
);
modport slave(
	input store,
	input store_idx,
	input store_data,
	output data
);

endinterface
