/*
 * Copyright (c) 2023 Robert Drehmel
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
module mmr_trigger_interface_connect(
	mmr_trigger_interface.master m,
	mmr_trigger_interface.slave s
);

for (genvar i = 0; i < m.N; i++) begin
	assign m.tsr_invpulses[i] = s.tsr_invpulses[i];
	assign s.tsr[i] = m.tsr[i];
end

endmodule
