/*
 * Copyright (c) 2023 Robert Drehmel
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */
module fifo_write_interface_connect(
	fifo_write_interface.master m,
	fifo_write_interface.slave s
);

assign m.clock = s.clock;
assign m.reset = s.reset;
assign m.wr_data = s.wr_data;
assign m.wr_en = s.wr_en;
assign s.full = m.full;
assign s.almost_full = m.almost_full;
assign s.wr_data_count = m.wr_data_count;

endmodule
